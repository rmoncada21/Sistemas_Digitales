// Circuito del ejercicio 4.1 modelado por comportamiento

module circuito (A, B, C, D, F1, F2)
    input A, B, C, D;
    output F1, F2;

    
endmodule